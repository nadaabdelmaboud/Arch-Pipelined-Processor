LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY MuxSignals IS
  PORT (
    IR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    ControlSignals : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
    CONTROL_HAZARD : IN STD_LOGIC;
    DATA_HAZARD : IN STD_LOGIC;
    OutSignals : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    OpCode : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END MuxSignals;

ARCHITECTURE a_MuxSignals OF MuxSignals IS
BEGIN

  OutSignals(13 DOWNTO 0) <= (OTHERS => '0') WHEN CONTROL_HAZARD = '1' OR DATA_HAZARD = '1'
ELSE
  ControlSignals(13 DOWNTO 0);

  OpCode <= (OTHERS => '0') WHEN CONTROL_HAZARD = '1' OR DATA_HAZARD = '1'
    ELSE
    IR(31 DOWNTO 26);
END a_MuxSignals;